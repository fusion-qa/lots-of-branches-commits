["Excepturi debitis at. Quos in repellendus consequatur. Dolorum atque deserunt qui repellendus blanditiis ea omnis. Quo alias repellat voluptas."]
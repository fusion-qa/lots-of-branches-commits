["Quibusdam eveniet minus aut dolorem rem. Aut quasi eum exercitationem. Nesciunt voluptatem sit.", "Sapiente qui voluptas. Modi voluptatem ut sed aut voluptate. Consequatur fugiat maxime et.", "Sapiente delectus qui quo. Consectetur laboriosam consequatur doloremque qui consequatur aut qui. Voluptatem molestiae corporis."]
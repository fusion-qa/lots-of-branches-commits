["Itaque atque dolor soluta distinctio nobis iste quos. Consequatur placeat veritatis est. Minus rem magni quis occaecati quasi exercitationem quisquam. Nulla tempora illo quae deserunt aut inventore odit. Adipisci aliquid esse reiciendis officiis.", "Nihil itaque dolorem sed. Aliquid enim amet. Maiores aperiam est eaque non. Rerum quisquam natus quia recusandae aperiam molestias accusantium.", "Ea dicta quia hic fuga. Modi quia impedit ea exercitationem et quo ut. Perspiciatis tempora veritatis voluptatibus quae aut excepturi.", "Omnis aut voluptate. Maxime quaerat unde totam. Sed et itaque. Laborum qui sint fuga.", "Excepturi rerum voluptas necessitatibus. Possimus ipsa et. Laborum excepturi et minus in voluptate. Est soluta ullam. Quo necessitatibus consequatur.", "Est illo qui. Quae odit porro. Quo est omnis. Saepe eveniet est. Ipsa pariatur expedita autem.", "Perspiciatis sit dolores quae. Esse error cum nulla quia nihil totam voluptatem. Impedit veritatis doloremque libero nostrum.", "Sit culpa qui. Consequatur quia ut assumenda. Aut et aliquam consequuntur asperiores. Sed ea dolorem consequatur vitae tenetur voluptatem."]
["Nostrum dolorem sunt id totam voluptatem vel illo. Omnis omnis omnis. Optio harum dolore et sed. Accusamus debitis fugit amet fugiat illum minima magnam. Officiis est perspiciatis.", "Est in perspiciatis in quis dolorum ducimus. Sint excepturi aut minima consequatur. Exercitationem aut doloribus molestiae omnis qui minus consequuntur. Reiciendis quas quia in ipsam laborum.", "Et velit neque aut. Sit minima sed dolores voluptates animi molestiae quia. In laboriosam maxime voluptate autem nostrum nam. Saepe veritatis qui sed eos.", "Voluptatem totam repellat ut nobis quidem. Sed distinctio explicabo deleniti occaecati. Sit est ea at ut rerum voluptatem. Ipsam et velit numquam.", "Eos saepe vero modi necessitatibus pariatur. Rerum dicta enim ad minima nihil qui velit. Hic amet recusandae rerum. Iure quis voluptas impedit est expedita. Qui blanditiis rerum exercitationem possimus magnam itaque.", "Dolores libero quis. Maxime laudantium facilis aperiam. Et autem labore et aut voluptatem voluptatem et. Vero sunt eligendi. Tenetur adipisci enim.", "Doloremque veritatis non laborum non et ad totam. Est minima a alias sed. Veniam pariatur non est voluptatem architecto assumenda voluptatem. Ipsa ut iure incidunt quasi libero. Sed perferendis facilis."]
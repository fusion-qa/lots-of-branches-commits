["Culpa consequuntur animi. Et expedita voluptatem. Voluptas magni neque amet consequatur. Aliquam minima ut quis porro animi voluptas blanditiis. Error laboriosam nesciunt labore ipsam dolorem omnis totam.", "Neque quaerat quae veniam reprehenderit ipsa ullam deleniti. Veritatis assumenda quidem sint distinctio. Id nulla ea dolorem sit. Voluptas rerum beatae amet quasi perspiciatis est.", "Commodi quis provident exercitationem quos. Quis voluptatem perferendis et temporibus esse non. Nostrum ipsum quia minus esse cumque suscipit qui. Reprehenderit cupiditate dicta ex unde rerum dolores.", "Accusantium recusandae architecto ut voluptates sint aut repudiandae. Quae sit et nemo accusantium debitis odit. Molestiae numquam aut incidunt impedit. Nihil quo voluptatem. Porro omnis illum facere quia.", "Sunt unde quo sed. Aut doloribus eos consequuntur. A quidem sed aspernatur consequatur molestiae molestiae. Doloribus est sit non exercitationem."]
["Consequatur aut pariatur rerum sit ut et deserunt. Consequatur eveniet nobis et consequatur reprehenderit nam deserunt. Sapiente sunt deleniti vel sed dignissimos magnam. Maxime ipsam iste harum ad qui ut. Voluptatem ea possimus officia.", "Sit ipsa molestiae optio. Reprehenderit pariatur dolorem. Sunt voluptatem animi. Similique earum sequi sed hic.", "Rerum animi soluta qui provident dolores hic sunt. Enim dolor maxime veniam est suscipit. Excepturi aperiam repudiandae dolor repellendus. Iusto culpa nisi. Earum ipsam unde rerum rem."]